----------------------------------------------------------------------------------
--                                LIBRARIES                                     --
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

----------------------------------------------------------------------------------
--                                 PACKAGE                                      --
----------------------------------------------------------------------------------

package serial_port_receiver_fsm_pkg is

  --------------------------------------------------------------------
  --                          COMPONENT                             --
  --------------------------------------------------------------------
  
  -- serial connection of flip-flops to avoid latching of metastable inputs at
  -- the analog/digital interface
  component serial_port_receiver_fsm is
    generic
    (
      CLK_DIVISOR : integer
    );
    port
    (
    clk, res_n, rx : in  std_logic;
    data_new : out std_logic;
    data                     : out  std_logic_vector(7 downto 0)
    );
  end component serial_port_receiver_fsm;
end package serial_port_receiver_fsm_pkg;
