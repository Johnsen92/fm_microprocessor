library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.pipeline_package.all;

package program_package is
    
    --constant MAX_PC : integer := 16; -- TODO: incl or excl, what is at last pc if anything
    constant MAX_PC : integer := 15;
    
    subtype PC_T is integer range 0 to MAX_PC;
    type INSTR_ARRAY_T is array(0 to MAX_PC) of INSTR_T;
--    constant PROGRAM : INSTR_ARRAY_T := (
--		"0101000000100011111111",
--		"0111010000100000001000",
--		"0110110000100011111111",
--		"0101000001000000000000",
--		"0101000001100000000000",
--		"0101000010000000000000",
--		"0101000010100000010010",
--		"0111010010100000001000",
--		"0110110010100001000111",
--		"0101000011000000000000",
--		"0101000011100001101101",
--		"0111010011100000001000",
--		"0110110011100011100000",
--		"0101000100000000001010",
--		"0001000100100111000000",
--		"0011000100100001000000",
--		"0001110100100000000000",
--		"0000110011000000000000",
--		"0010010011000000000000",
--		"0001010001000101000000",
--		"0001000011000010000000",
--		"0010000011100010000000",
--		"1001100000000000011000",
--		"0001000001001001000000",
--		"1111110100000000000000",
--		"1000000000000000010001",
--		"0000000000000000000000"
--    );
    
    constant PROGRAM : INSTR_ARRAY_T := (
        OP_MOVI & "00001" & "00011111111",               --1: 0000001001001001
		OP_SLL	& "00001" & "00000001000",
		OP_MOVI	& "00010" & "00011010101",
		OP_SLL	& "00010" & "00000001000",
		OP_SUB	& ""
        (others => '0')
    );

end program_package;