PACKAGE sp_const_pkg IS
	CONSTANT DATA_WIDTH : INTEGER := 8;
	CONSTANT BAUD_RATE : INTEGER := 115200;
	CONSTANT TX_FIFO_DEPTH : INTEGER := 10;
	CONSTANT RX_FIFO_DEPTH : INTEGER := 10;
	CONSTANT CLK_FREQ : INTEGER := 25000000;
END PACKAGE sp_const_pkg;
